﻿return {

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_import = "Ett fel uppstog vid importering av tilläggsmodul.",
    msg_usage = "Användning: [+!#]unban ip|nick|cid <IP>|<ANVÄNDARNAMN>|<CID>",
    msg_off = "Hittade inte användaren.",
    msg_god =  "Du har inte behörighet att ta bort användarens bann.",
    msg_ok = "Användare %s tog bort bannen på %s.",

    help_title = "cmd_unban.lua",
    help_usage = "[+!#]unban ip|nick|cid <IP>|<ANVÄNDARNAMN>|<CID>",
    help_desc = "Unbannar användare efter IP, ANVÄNDARNAMN eller CID",

    ucmd_menu_ct1_1 = { "Användare", "Kontroll", "Unban", "efter NICK" },
    ucmd_menu_ct1_2 = { "Användare", "Kontroll", "Unban", "efter CID" },
    ucmd_menu_ct1_3 = { "Användare", "Kontroll", "Unban", "efter IP" },

    ucmd_ip = "IP-adress:",
    ucmd_cid = "CID:",
    ucmd_nick = "ANVÄNDARNAMN:",

}