﻿return {

    client_mode_a = "aktiv",
    client_mode_p = "passiv",
    client_ssl_n = "nej ( aktivera gärna det! )",
    client_ssl_y = "ja",

    msg_ccpm_1 = "ja ( aktiverat för din åtkomstnivå )",
    msg_ccpm_2 = "ja ( inaktiverat för din åtkomstnivå )",
    msg_ccpm_3 = "nej",

    msg_years = " år, ",
    msg_days = " dagar, ",
    msg_hours = " timmar, ",
    msg_minutes = " min, ",
    msg_seconds = " sek",

    msg_unknown = "<OKÄNT>",

    msg_info_1 = [[


=== ANVÄNDARENS INLOGGNINGSINFO ==============================

        Användarnamn:	%s
        IP-adress:	%s
        Åtkomstnivå:	%s  [ %s ]

        Klientversion:	%s
        Klientläge:	%s
        Klient-SSL:	%s
        Klient-CCPM:   %s

        Registrerad av:	%s
        Registrerad den:	%s

        Senast inloggad:  %s

        TLS-läge:   %s
        TLS-cipher:  %s

============================== ANVÄNDARENS INLOGGNINGSINFO ===
   ]],


    msg_info_2 = [[


=== ANVÄNDARENS INLOGGNINGSINFO ==============================

        Användarnamn:	%s
        IP-adress:	%s
        Åtkomstnivå:	%s  [ %s ]

        Klientversion:	%s
        Klientläge:	%s
        Klient-SSL:	%s
        Klient-CCPM:   %s

        Registrerad av:	%s
        Registrerad den:	%s

        Senast inloggad:  %s

        TLS-läge:   %s
        TLS-cipher:  %s

        Hubbversion:	%s

============================== ANVÄNDARENS INLOGGNINGSINFO ===
   ]],

}