﻿return {

    help_title = "cmd_restart.lua",
    help_usage = "[+!#]restart [<MEDDELANDE>]",
    help_desc = "Startar om hubben",

    ucmd_menu = { "Hubb", "Kärna", "Omstart av hubben", "KLICK" },
    ucmd_msg = "Gruppmeddelande (valfritt)",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_ok = "Hubben startar om...",

    msg_countdown = "*** Omstart av hubben om ***",

    msg_restart = [[


=== OMSTART AV HUBBEN ======================================================================================================

  %s

====================================================================================================== OMSTART AV HUBBEN ===

  ]],

}