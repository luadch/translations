﻿return {

    client_mode_a = "aktiv",
    client_mode_p = "passiv",
    client_ssl_n = "nej ( aktivera gärna det! )",
    client_ssl_y = "ja",

    msg_ccpm_1 = "ja ( aktiverat för din åtkomstnivå )",
    msg_ccpm_2 = "ja ( inaktiverat för din åtkomstnivå )",
    msg_ccpm_3 = "nej",

    msg_years = " år, ",
    msg_days = " dagar, ",
    msg_hours = " timmar, ",
    msg_minutes = " min, ",
    msg_seconds = " sek",

    msg_unknown = "<OKÄNT>",

    msg_info = [[


=== ANVÄNDARENS INLOGGNINGSINFO ==============================

        Användarnamn:	%s
        IP-adress:	%s
        Åtkomstnivå:	%s  [ %s ]

        Klientversion:	%s
        Klientläge:	%s

        Registrerad av:	%s
        Registrerad den:	%s

        Senast inloggad:  %s

        Klient-SSL:	%s
        TLS-läge:	%s
        TLS-cipher:	%s

============================== ANVÄNDARENS INLOGGNINGSINFO ===
   ]],

}