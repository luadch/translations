﻿return {

    help_title = "cmd_rules.lua",
    help_usage = "[+!#]rules",
    help_desc = "Visar hubbens regler",

    ucmd_menu =  { "Allmänt", "Regler" },

}