﻿return {

    help_title = "etc_cmdlog.lua",
    help_usage = "[+!#]cmdlog show",
    help_desc = "Visar kommandologgen",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_nofile = "Hittade ingen 'cmd.log'",
    msg_usage = "Användning: [+!#]cmdlog show",

    msg1 = "   |   Kommando: [+!#]",
    msg2 = "   |   använd av: ",

    msg_out = [[

    
=== KOMMANDOLOGGARE ========================================================================================

%s
======================================================================================== KOMMANDOLOGGARE ===

      ]],

    ucmd_menu = { "Hubb", "Loggar", "visa", "cmd.log" },

}