﻿return {

    client_mode_a = "M:A ( aktiv )",
    client_mode_p = "M:P ( passiv )",
    client_ssl_n = "NEJ ( aktivera gärna det! )",
    client_ssl_y = "JA",

    msg_ccpm_1 = "JA ( aktiverat för din åtkomstnivå )",
    msg_ccpm_2 = "JA ( inaktiverat för din åtkomstnivå )",
    msg_ccpm_3 = "NEJ",
    
    msg_days = " dagar, ",
    msg_hours = " timmar, ",
    msg_minutes = " min, ",
    msg_seconds = " sek",
    
    msg_unknown = "<okänt>",

    msg_info_1 = [[


=== ANVÄNDARENS INLOGGNINGSINFO =======================

        Användarnamn:	%s
        IP-adress:	%s
        Åtkomstnivå:	%s  [ %s ]

        Klientversion:	%s
        Klientläge:	%s
        Klient-SSL:	%s
        Klient-CCPM:   %s

        Registrerad av:	%s
        Registrerad den:	%s
        
        Senast inloggad:  %s

======================= ANVÄNDARENS INLOGGNINGSINFO ===
   ]],


    msg_info_2 = [[


=== ANVÄNDARENS INLOGGNINGSINFO =======================

        Användarnamn:	%s
        IP-adress:	%s
        Åtkomstnivå:	%s  [ %s ]

        Klientversion:	%s
        Klientläge:	%s
        Klient-SSL:	%s
        Klient-CCPM:   %s

        Registrerad av:	%s
        Registrerad den:	%s
        
        Senast inloggad:  %s


        Hubbversion:	%s

======================= ANVÄNDARENS INLOGGNINGSINFO ===
   ]],

}