﻿return {

    help_title = "cmd_errors.lua",
    help_usage = "[+!#]errors",
    help_desc = "Visar error.log",

    ucmd_menu =  { "Hubb", "Loggar", "visa", "error.log" },

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_noerrors = "Inga fel",

}