﻿return {

    help_title = "cmd_slots.lua",
    help_usage = "[+!#]slots",
    help_desc = "Visar användare med lediga slottar",

    ucmd_menu =  { "Användare", "Lediga slottar" },
    
    msg_out = [[


=== LEDIGA SLOTTAR ====================

%s
==================== LEDIGA SLOTTAR ===
  ]],

}