﻿return {

    msg_banner = [[


    === BANNER ================================================================

                ::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::
                :::::::::::::::::   ::::::::::::::::::::::::::::::::::::::::::::::::::::::   ::::::::::::::::::   ::::::::::::::::::::::::::::::
                :::::::::::::::::    :::::::::::::::::::::::::::::::::::::::::::::::::::::    :::::::::::::::::    :::::::::::::::::::::::::::::
                :::::::::::::::::    :::::::::::::::::::::::::::::::::::::::::::::::::::::    :::::::::::::::::    :::::::::::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   ::::            ::::::            :::::          ::            :::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   ::::             ::::             ::::          :::             ::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   ::::::::::::::   :::    ::::::    :::    ::::::::::    :::::    ::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   ::::::           :::   :::::::    ::    :::::::::::    ::::::   ::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   ::::             :::   :::::::    ::    :::::::::::    ::::::   ::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   ::::             :::   :::::::    ::    :::::::::::    ::::::   ::::::::::::::::::::
                :::::::::::::::::    ::::::::::    ::::::   :::    :::::::   :::   :::::::    ::    :::::::::::    ::::::   ::::::::::::::::::::
                ::::::::::::::::::     :::::::::    :::::   :::    :::::::   :::     :::::    :::     :::::::::    ::::::   ::::::::::::::::::::
                :::::::::::::::::::           ::            ::::             ::::             ::::           ::    ::::::   ::::::::::::::::::::
                :::::::::::::::::::::         ::::          :::::            ::::::          ::::::         :::   :::::::   ::::::::::::::::::::
                ::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::
                Luadch hemsida: http://luadch.github.io

    ================================================================ BANNER ===
      ]],

}