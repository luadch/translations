﻿return {

    msg_sharelimits = "Minsta/högsta utdelning i hubben: %s/%s  Din utdelning: %s",

}