﻿return {

    msg_denied = "Du har inte behörighet att använda detta kommando eller så har användare högre åtkomstnivå än dig.",
    msg_usage = "Användning: [+!#]upgrade sid|nick|cid <SID>|<ANVÄNDARNAMN>|<CID> <ÅTKOMSTNIVÅ>",
    msg_off = "Hittade inte användaren.",
    msg_reg = "Användaren är inte registrerad eller så är det en bot.",
    msg_out = "%s  ändrade  %s  från åtkomstnivå: %s [ %s ]  till:  %s [ %s ]",
    msg_out_2 = "%s  med åtkomstnivå:  %s [ %s ]  har försökt ändra  %s  till:  %s [ %s ]",
    msg_same = "Användaren har redan denna åtkomsnivå, inga ändringar behöver göras.",

    help_title = "cmd_upgrade.lua",
    help_usage = "[+!#]upgrade sid|nick|cid <SID>|<ANVÄNDARNAMN>|<CID> <ÅTKOMSTNIVÅ>",
    help_desc = "Ställer åtkomstnivå på användaren",

    ucmd_menu = "Uppgradera",
    ucmd_level = "Åtkomstnivå:",
    ucmd_popup = "Använarnamn:",
    
    ucmd_menu_ct1_1 = "Användare",
    ucmd_menu_ct1_2 = "Kontroll",
    ucmd_menu_ct1_3 = "Uppgradera",
    ucmd_menu_ct1_4 = "efter ANVÄNDARNAMN från lista",
    ucmd_menu_ct1_5 = "Användare",
    ucmd_menu_ct1_6 = "Kontroll",
    ucmd_menu_ct1_7 = "Uppgradera",
    ucmd_menu_ct1_8 = "efter ANVÄNDARNAMN",

}