﻿return {

    help_title = "cmd_restart.lua",
    help_usage = "[+!#]restart [<MEDDELANDE>]",
    help_desc = "Startar om hubben",

    ucmd_menu = { "Hubb", "Kärna", "Hubbomstart", "KLICK" },
    ucmd_msg = "Gruppmeddelande (valfritt)",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_ok = "Hubbomstart...",

    msg_countdown = "*** Omstart av hubben om ***",

    msg_restart = [[


=== HUBBOMSTART ======================================================================================================

  %s

====================================================================================================== HUBBOMSTART ===

  ]],

}