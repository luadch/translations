﻿local lang = {}
lang.pics = {}

lang.help_title = "cmd_ascii.lua"
lang.help_usage = "[+!#]ascii <NAMN>"
lang.help_desc = "Visar en <ASCII-BILD> i huvudchatten; Lista över alla bilderna: "
lang.help_err = "Kunde inte hitta bilden"

lang.ucmd_menu =  { "Allmänt", "Ascii" }

lang.pics.afk = function(user) return [[



             ()::()    
          (´( 'o' )    
           ,-(___)_'--.   
       =(o)===(o)='

 ]]..user..[[ är inte här...


	]]
end

lang.pics.lol = function(user) return [[



 	           ,.·^*''l'\            .·^*'´¯¯¯''*^·,.  ,/l''*^·-,
 	           'l       'l::\       ,·'     ,.·:*:·,     ''i::; 'l          l
 	           'l       'l:::      ;       ':,:::,:·       ';:::'l          l'
 	           'l       l::;i - ·;i' :,      ¯¯       ,·´l::::'l          l
 	           'l       '´       'l'i::: *: ·.–·    ^*'´: :'l::,.       '''*· ,
 	           'l        ,.-:^:':'\:' :;:: :: : : : :: ::; ·'i:::l':^·.,     ''i
 	           'l  ,.:'':::::::::::'\  ' *^ ·:–:· ^*'´  'l/::::::::''::^:. ,l
 	           '´:;:::::::::;:-·^*'                             '*^·:;-L:;·'
 	               '·;:·'                                               '^·:;·''


	]]
end

lang.pics.hej = function(user) return [[



            ,;'’¨¯'·¸ ¸.· ;'''ˆ’¨¯¯ˆ¯’¨¨;.,;'’¨¯'·¸
            'l        .´_ .    ¨¨ .,,,·    ¹ ¹         l
             `'-,,    ;,¨o¨ ¸   ¸.´ o  ';   '.¸    ,--'
                  '  ;  .¸,.-˜   '·.¸_¸·       ˜;'
                   -˜    ¸˜ I ˜·¸   ¸          ¸'
                   `-,    ' -^- -'         ¸ ¸.·'
                       ¸'  --...,- -     `'l
                    ,  :;´´              `**-;,
   -------------ooOOo-------oOOoo----------------------------

         Hej :D
         ]]..user..[[  det är dags för lite småprat :D


	]]
end

lang.pics.hej2 = function(user) return [[



 		                                    oooooooooooooooooooo
 		                              oo0000000000000000000000o
 		                          oo000000000000000000000000000o              o0   00   o0
 		      o 0  oo      o000000000000000000000000000000000o       00 00  00o
 		oo  0 0  0      o000000000      0000000000       000000000o         000o00o0
 		 000000o0    o000000000   #     000000000  #   0000000000o      0000000
 		  0000000   00000000000        000000000         00000000000000000000000
 		  000000000000000000000    00000000000     0000000000000        000
 		    000    00000000000000000000000000000000000000000000          000
 		    000    o000000000000000000000000000000000000000000000          000o
 		   o00    00000000000000000000000000000000000000000000000           000o
 		   000    0000000000000000000000000000000000000000    0000000ooooo0000o
 		  o000oo00000  0000000000000000000000000000000000    o000 0000000000000
 		  000000 0000   000000000000000000000000000000000   0000
 		              0000     000000000000000000000000000000          o000
 		                000o        00000000000000000000000000           0000
 		                 000o                     0000000000000000                 o000
 		                  0000o         ****** BÄÄÄÄÄÄÄÄÄÄH******    o000
 		                    0000o          o0000000o 0000000o           o0000
 		                     00000oo       0000000o00000000o    o0000
 		                         0000ooo     0000000o0000000000000
 		                            000000oo   00000000000000000
 		                                           000000000000000000
 		                                            000000000000000000.
 		                                              00000000000000000
 		                                                  0000000000000

 BOOOOOH
 ]]..user..[[ är här...


	]]
end

lang.pics.hej3 = function(user) return [[



            ;::::; :;
          ;:::::'   :;
         ;:::::;     ;.
        ,:::::'       ;           OOO
        ::::::;       ;          OOOOO
        ;:::::;       ;         OOOOOOO
       ,;::::::;     ;'         * OOOOOOO
     ;::::::::: . ,,,;.        *  * DOOOOO
   .';:::::::::::::::::;,     *  *     DOOOO
  ,::::::;::::::;;;;::::;,   *  *        DOOO
 ; :::::: '::::::;;;::::: ,#*  *          DOOO
 : ::::::: ;::::::;;::: ;::#  *            DOOO
 :: ::::::: ;:::::::: ;::::# *              DOO
  : ::::::: ;:::::: ;::::::##               DOO
  ::: ::::::: ;; ;:::::::::##                OO
  :::: ::::::: ;::::::::;:::#                OO
   ::::: ::::::::::::;' :;::#                O
    ::::: ::::::::;' *  *  :#
    :::::: :::::;'  *  *    #

 Den obarmhärtigt själsökaren ]]..user..[[ är här...


	]]
end

lang.pics.morgon = function(user) return [[



 ___ ___
I     V     I
I       ORNING
I__IVI__I
 __    __
I    I_I    I
I     _  AVE A NICE
I__I  I__I
 ___
I       ' .
I    D   i
I.___, 'AY

 ]]..user..[[  önskar er en god morgon !


	]]
end

lang.pics.morgon2 = function(user) return [[



   ,XX    ,§§,    ,;;;,
  (  ö, )  ( ü  )  (  ö )
   (') (')   (') (')   (') (')

 Dessa 3 & ]]..user..[[ önskar dig en stressfri, motiverande dag!


	]]
end

lang.pics.sova = function(user) return [[



 ---------  --------------------------------------------------------------------------------------------
 ---------
 ---------
 ---------                                           zzz
 ---------                                               ZZZ
 ---------                                                       zz
 ---------     o                                                    zz    _ .-----.      ___ O
 ---------     l l                                                         )          `. ,'         l l     
 ---------     l l                                                     (` '               l        : l         trevliga
 ---------     l l                                     _..-.-.-.-._    )       , )     ,'.        l l                drömmar...
 ---------     l l ( ' .                     __..- '    ) ) ) ) ) )``-'               . -          l l  
 ---------     l l    `...------''``--'''''    )_______....---      _, -- ' '                 ; l
 ---------     l l__(_..-......____..._,-'_,..____....__..- '  ..________ ..' l l
 ---------     l l_________________________________________l l
 --------- __l_l________________________________________l_l__
 ---------

            ]]..user..[[  går och lägger sig...


	]]
end

lang.pics.sova2 = function(user) return [[



 			                                 ___       .
 			 .    *                  _.--'   __'-.
 			                      ,-'        .-      '-\
 			                      ,-'        .-      '-\              .
 			     *   .          .^         /           ( )      .
 			              +   {_.---._/
 			                   /      .  Y
 			        *        /        \_j         *             +
 			   .             Y     ( ool__            ***Godnatt hubbsters***
 			                _             '-.           .
 			                _      (___      \
 			         .      _        .)   -.__/             .
 			                 l        _)
 			 .                 \      'l              *
 			     +              \       ^.
 			                        '-._       -.___,
 			                   .         '--..____.^
 			*                                 .                      *

            ]]..user..[[  går och lägger sig...


	]]
end

lang.pics.sova3 = function(user) return [[



                                                 ·´`·.(*·.¸(`·.¸ ¸.·´)¸.·*).·´`·
                                    ·´¨*·.¸¸          GODNATT         .¸¸.·*¨`·
                                                 ·´`·.(¸.·´(¸.·* *·.¸)`·.¸).·´`·

                                     ]]..user..[[  går och lägger sig...


	]]
end

lang.pics.sova4 = function(user) return [[



                         boing         boing         boing
               e-e           . - .         . - .         . - .
              (\_/)\       '       `.   ,'       `.   ,'       .
               `-'\ `--.___,         . .           . .          .
                  '\( ,_.-'
                     \\               ``             ``
                     ^'          Hoppar in i drömlandet...   Godnatt...

                  ]]..user..[[  går och lägger sig...


	]]
end

lang.pics.sova5 = function(user) return [[



    *      +    *      *   +     *
    *   + *  God     *  +    *
   +     *  +  Natt *  +  *   +    *
   +    *  +   *      +   *   +   +
     +*   *   +   *   * +   + +   + +
    *   *  +  ]]..user..[[ *   +
    + + **  +  går till sängs * +   *
      +      *    + *    +   +  *  + *


	]]
end

lang.pics.thc = function(user) return [[



                                   .:.
                                   :_:
                                  .:_:.
                                  ::_::
                   :.             ::_::             .:
                   :_:.          .::_::.          .:_:
                   ::_:.         :::_:::         .:_:;
                    ::_:.        :::_:::        .:_::'
                    ::_::.       :::_:::       .::_:;
                     ::_::.      :::_:::      .::_::'
                     :::_::.     :::_:::     .::_::;
                      :::_::.    :::_:::    .::_::;'
             ::.       :::_::.   :::_:::   .::_::;'      .:;'
              :::..     :::_::.  :::_:::  .::_::;'    ..::;'
               ::::::.   :::_::. :::_::: .::_::;'  .:::::;'
                  ::::::. :::_::.:::_::;.::_::;'.:::::;'
                    ::::::. ::_::.::_::.::_::'.:::::;'
                       :::::::::_:::_:::_::::::::;'
                           :::::::_:_::_:::::;''
                               ::::::::::;'
                             .:;'' :::   ::.
                                  : : :

                   ]]..user..[[ är stenad !


	]]
end

lang.pics.thc2 = function(user) return [[



 		           ;::::;
 		           ;::::; :;
 		         ;:::::'   :;                                      ( ( (  )
 		        ;:::::;     ;.                                    ( ) ( ´)
 		       ,:::::'  00 ;                                  ( ( ' )
 		       ::::::;   J_______,.,.,.,.___l    ( (
 		       ;:::::;   (_______l l l l l____] '
 		      ,;::::::;     ;'          *¨¨¨¨¨´*
 		    ;::::::::: . ,,,;.        l  *  * /
 		  .';:::::::::::::::::;,     l      /
 		 ,::::::;::::::;;;;::::;,   l  *  /
 		; :::::: '::::::;;;::::: ,#*  /
 		: ::::::: ;::::::;;::: ;::#  *
 		:: ::::::: ;:::::::: ;::::# *
 		 : ::::::: ;:::::: ;::::::##
 		 ::: ::::::: ;; ;:::::::::##
 		 :::: ::::::: ;::::::::;:::#
 		  ::::: ::::::::::::;' :;::#
 		   ::::: ::::::::;' *  *  :#
 		   :::::: :::::;'  *  *    #

           Wow, det smakar bra, ]]..user..[[  rökar det finaste gräset i stan :D


	]]
end

lang.pics.beer = function(user) return [[



                    o*O8*.o..
           _o8O0o0OoO8OO.
          I         .    .    .      '80
  .===[I         :    ;    :      Io°O
 II       I        :    ;   :        I°o
 II       I        :    ;   :        I°
 II       I        :    ;   :        I
 II       I        :    ;   :        I
  '===[I         .    .    .      I
          I_____________I


   ]]..user..[[ : det är dags för en kall öl :D


	]]
end

lang.pics.cigg = function(user) return [[



     ( (
      ) )    Det är dags för en cigarett  !
     ( (
       ___________________
      ()_______________)::)::)

 ]]..user..[[ röker...


	]]
end

lang.pics.nodispute = function(user) return [[



                 ()()
                (._.)
             (')(')_)

     No Dispute! otherwise I come!


	]]
end

lang.pics.kaffe = function(user) return [[



 			                )
 			              ( (             Kaffedags
 			           (`````)o
 			          '''''''''''''

             ]]..user..[[  dricker en kopp...


	]]
end

lang.pics.bad = function(user) return [[



                 o      .   _       .
                    .       (_)           o
       o             ____                         _         o
      _          ,-/        /)))        .     o  (_)   .
     (_)        \_\   ( e e)          O            _
  o                 \  / '  _/     ,_ ,  o    o    (_)
    .   O         _/    (_      / _/       .   ,           o
            o8o/           \_ / /  .,-.,       oO8    / ) 
      o8o8O l       }   } /  /   \Oo8OOo8Oo  l  l     O
        Oo (''''''o8'''''''''''''''''''''''''''''''''''''''''''''''''8oo'''''''''''''''''')
      _       \`'                                                `'   /'   o
     (_)       \                                                     /     _   .
          O      \                                                 /     (_)
    o         .    \_______________________/
              --------(_/----------------------------\_)--------

 ]]..user..[[ hoppar snabbt i badet...


	]]
end

lang.pics.telefon = function(user) return [[



            _______
      @ (_)---------(_)
   @      /  ### \    *RING*
   @     /   ###  \     *RING*
  @ @/    ###    \
          ¯¯¯¯¯¯¯¯¯

 ]]..user..[[  ringer...


	]]
end

lang.pics.omstart = function(user) return [[



                          o
                          I        o
                          I    o   I
                          I    I    I
                  l'''''''''''''''''''''''''''''''''''''l
             l''''''''''''''''''''''''''''''''''''''''''''''''''''l
        l''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''l
  l''''''''''''''''       OMSTART       ''''''''''''''''l
  ''''''''l_______________________l''''''''
             l_________________l
                     /                \
                     ''''''''''''''''''''''''''''''
                        *      *     *
                   *    *    *       *    *
               *    *    *       *    *  *    *

 ]]..user..[[  måste starta om sin fickkalculator :D


	]]
end

lang.pics.sjuk = function(user) return [[



     o>
i , /(,_,
I==========I
Jag är sjuk!

i ,o_,__,
I==========I
Jag måste gå och lägga mig...")

 ]]..user..[[  är sjuk :-o


	]]
end

lang.pics.leakme = function(user) return [[



  	      ¸.-•˜˜˜˜¨¨˜_•.¸
 	       ¸˜¸,.¸    ¸,..¸  ˜¸
 	       _¸o›¸ ‹ o›  __¸˜.,,¸¸___
 	       (¸ (_,     )¸/˜¸;;;;;;;;;;;;;;˜•-.,¸
 	        ¨˜\,¸.´_ ¸--- ¸  ;;;;;;;;;;;;;;;;;;;;;¸
 	         (_¸.•¸˜;;;;;;;¸;;;;;;;;;;;;;;;;;;;;;;;;;;-,¸ 
 	               ˜¸;;;;;;; _¸ ;;;;;;;;;;;;;;¸¸¸.••-••˜˜˜˜˜•-.¸
 	                  ˜¸.•˜˜˜ ¸;;;;;;;;˜¸•˜          •¸         ˜•¸
 	                    ˜¸     ˜¸';;;¸,¸˜               ˜¸         ˜¸
 	                       ˜,   ˜¸;;;;;_                  _         _
 	                         ˜¸   \¯¯˜¸                 _        ¸˜¸
 	                           ˜¸  ˜¸ ¸-˜¸¸¸,,..---••••••˜˜˜˜˜˜˜¨¨¨¯•¸
 	                           ¸˜ ,¸  ¸˜•••••˜˜¨¨•••:::::::::::::::••˜¨¸˜
 	                            ˜• ¸_ ˜¸      ¸ ¯;¸ ´ ¸-•¨  ¸ ¯¸ ´  ¸˜
 	                                ¯¯ ˜¸   _¨˜˜¨     ¯¸   ¨˜˜¨      ˜¸
 	                                     ˜•¸   •˜¸--¯  ˜•.¸ •˜¸-•-•¸¨ ˜¸
 	                                        '¸      ¯      \¸          ˜¸
 	                                       ¸.˜__,..-..¸-•˜__,..-.,,_\¸
 	                                      (;;;;;;;;˜;;;;;¸\¯\¸;;;;;;;;;)˜˜

  Leak me!  *gg*
  ]]..user..[[  låter tankarna flöda...


	]]
end

lang.pics.pask = function(user) return [[



          ***
         ** **
        **   **
        **   **         ****
        **   **       **   ****
        **  **       *   **   **
         **  *      *  **  ***  **
          **  *    *  **     **  
           ** **  ** **        **
           **   **  **
           *            *
        *                  *
      *      0       0      *
     *     /    @           *
      *    __/ __/        *
       *         W         *
          **           **
              *****

 Glad Påsk önskar ]]..user..[[ !


	]]
end

lang.pics.lyssna = function(user) return [[



       .²´¯¯¯¯¯'‚
           '' ,''.      '.
                   '.,  .;
                     ;  ;
                     ,. ,
                     '¸ ¸.· ;'''ˆ'¨¯¯ˆ¯'¨¨;·.,;'''¨¯'·¸
                     .´_ .    ¨¨ .,,,·    ¹  ¹        .¹
                    ;,¨o¨ ¸   ¸.´ o ';    '.¸         '¸
                   ';  .¸,.-˜   '·.¸_¸·        ˜·¸     '¸
              ¸.¸.-·˜      ¨¯¨     ¸,.-¸        ¸'     '¸
            ¸˜   ˜·¸             ¸·˜ ¸.·˜    ¸,.·˜'·.¸   ˜·¸
             ˜·.¸¸.˜            ¸˜ ¸'       ¸'          ˜·-..˜¸
                ˜¸,,.--..,¸,.-·˜¸.·˜    ¸.·
                         ¸´,.- '   ¸,·*'
                            ·-·-· ´

 ]]..user..[[ lyssnar uppmärksamt på...


	]]
end

lang.pics.glad = function(user) return [[



 	 ,;' .;:                         *    ..:
 	  ::.        ..:,:;.,:;.       ;;     ::     .::::.
 	   ```::,      ::  ::  ::     ::     ::    ;:   .::
 	 ,:`;  ::;    ::  ::  ::     ::     ::    ::,::``
 	  :,,,,;;`  ,;; ,;;, ;;,  ,;;,   ,;;,   :,,,,:`

  ]]..user..[[ finner allt mycket underhållande...


	]]
end

lang.pics.ros = function(user) return [[



     { --.-'_,}
   {; \,__.-'}
   {.'- .__;-';
     '--.__.-'
       .-\\,-''-.
        - \( '-. \
           \;---,/
      .-''''-;\
     /  .-' )\
     \,---'  \

 Stressa ej, var glad!
 Denna ros är en gåva från  ]]..user..[[


	]]
end

lang.pics.nyfiken = function(user) return [[



                                                      .-- '' ~~ ''  ~''\___
                                                    Y                    !  ~~''\
                                                     !    `v. , _    _/''          !
                                                     \     ]      7~~''         /'
                                                       \   ]    / / ~''------''~
                                                    __.} ]_/-^-<-.
                                             .--''~        Y       ]  Y
                                           /                ]      oj-<______
                                         Y            _     ~---~    (      ^  Y
                                          [            !~t-.__(     // \. _ . ^
                                           \          ! !      ~\         _.^
                                             ''-._    ! !          ''---''~
                                                  Y  !-^----------.., __
                     .                             !  !--.,__   --.,__  ~ ''-.
                      \\                          !  ! !    ''~--.,_  ~--.     \
                        \\       _____       !  \ \___ ,      ''-._     /
                          \>-''~         ~''-.--j    ~------ /          ''--''
                          /              , -- .               Y
                      _Y_ /           (     )      ___  ]_
                 ,-~   ''                 ''--''      ''   ~- <   ~ -.
               /                                Y              \        \
             /               /         .        ]                  Y   )  Y
           /          ]    / -.____[        ]\,            )  !   /  /
        Y       /  /''--''  /         \ __ /'   \         / /_K-~
        `\__K-'' \__.-''                         ^.__K-''

  VAD? VEM? VAR?
  ]]..user..[[ är nyfiken...


	]]
end

return lang