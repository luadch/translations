﻿return {

    msg_slotlimits = "[ ANVÄNDARSLOTTAR ]--> Minsta antalet slottar i hubben:  %s  |  Högsta antalet slottar i hubben:  %s  |  Dina slottar:  %s",
    msg_redirect = "[ ANVÄNDARSLOTTAR ]--> Du blev omdirigerad därför att:  ",

}