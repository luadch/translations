﻿return {

    msg_sharelimits = "[ ANVÄNDARUTDELNING ]--> Lägsta utdelningsgränsen i hubben:  %s  |  Högsta utdelningsgränsen i hubben:  %s  |  Din utdelning:  %s",
    msg_redirect = "[ ANVÄNDARUTDELNING ]--> Du omdirigerades eftersom:  ",

}