﻿return {

    help_title = "cmd_hubstats.lua",
    help_usage = "[+!#]hubstats",
    help_desc = "Visa statistik om hubben",

    ucmd_menu_ct1 = { "Hubb", "etc", "Hubbstatistik" },

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_empty_tbl = "\n\n\tDen första statistiken kommer att synas i slutet av nästa månad.\n",
    msg_label = "\tÅR\t\tMÅNAD\t\tØ ANVÄNDARE\tØ UTDELAT\tREGISTRERINGAR\t\tAVREGISTRERINGAR\tBAN's\t\tUNBAN's",
    msg_stats = [[


=== HUBBSTATISTIK ========================================================================================================================

%s
%s
%s
======================================================================================================================== HUBBSTATISTIK ===
  ]],

}