﻿return {

    msg_invalid = "Ogiltig namngiven parameter i inf: ",

}