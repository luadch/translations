﻿return {

    help_title = "cmd_shutdown.lua",
    help_usage = "[+!#]shutdown",
    help_desc = "Stänger ner hubben",

    ucmd_menu = { "Hubb", "Kärna", "Hubbnerstängning", "KLICK" },

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_ok = "Stänger ner hubb...",

    msg_countdown = "*** Hubben stängs ner om ***",

}