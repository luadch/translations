return {

report_msg = "[ MISSLYCKAD INLOGGNING ]--> Användaren:  %s  |  IP:  %s  |  CID:  %s  |  Anledning:  %s",

}