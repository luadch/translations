﻿return {

    msg_sharelimits = "Minsta delning i hubben: %s  |  Max delning i hubben: %s  |  Din delning: %s",

}