﻿return {

    msg_denied = "Du har inte behörighet att använda denna chatten.",
    msg_send = "Ditt meddelande är skickat till alla Operatörer.",
    msg_toops = "Nytt %s meddelande från: %s | Msg: %s",

}