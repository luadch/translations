﻿return {

    help_title = "etc_topic.lua",
    help_usage = "[+!#]topic <NYTT_ÄMNE>",
    help_desc = "sätt hubbämne",

    msg_topic_changed = "%s har ändrat hubbämnet till: %s   |   det gamla hubbämnet var: %s",
    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_usage = "Användning: [+!#]topic <NYTT_ÄMNE>",

    ucmd_popup = "Nytt ämne:",
    ucmd_menu = { "Hubb", "Kärna", "Sätt hubbämne" },

}