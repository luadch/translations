﻿return {

    msg_denied = "[ TA BORT ]--> Du har inte behörighet att använda detta kommando eller att ta bort användarkonton med denna åtkomstnivå.",
    msg_usage = "Användning: [+!#]delreg nick <ANVÄNDARNAMN>  /  eller ta bort med svartlistspost:  [+!#]delreg nick <ANVÄNDARNAMN> <BESKRIVNING>",
    msg_error = "[ TA BORT ]--> Ett fel uppstod: ",
    msg_del = "[ TA BORT ]--> Ditt konto har tagits bort.",
    msg_bot = "[ TA BORT ]--> Användaren är en bot.",
    msg_ok = "[ TA BORT ]--> Användaren:  %s  har tagits bort av:  %s",
    msg_ok2 = "[ TA BORT ]--> Användaren:  %s  har tagits bort och svartlistad av:  %s  |  anledning: %s",
    msg_notfound = "[ TA BORT ]--> Användaren är inte registrerad.",

    help_title = "cmd_delreg.lua",
    help_usage = "[+!#]delreg nick <ANVÄNDARNAMN>  /  eller ta bort med svartlistspost:  [+!#]delreg nick <ANVÄNDARNAMN> <BESKRIVNING>",
    help_desc = "Ta bort en användare",

    ucmd_menu_ct1 = { "Användare", "Kontroll", "Delreg", "efter ANVÄNDARNAMN" },
    ucmd_menu_ct2 = { "Delreg", "OK" },
    ucmd_nick = "Användarnamn:",
    ucmd_reason = "Anledning: (läggs inte i svartlistan om den är tom)",

}