﻿return {

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_nochange = "Inga förändringar behövs.",
    msg_usage = "Användning: [+!#]setpass nick <ANVÄNDARNAMN> <LÖSENORD>  /  [+!#]setpass nick myself <LÖSENORD>",
    msg_god = "Du har inte behörighet att ändra lösenordet på denna användaren.",
    msg_reg = "Användaren är inte registrerad eller så är det en bot.",
    msg_ok = "Lösenordet har ändrats till: ",
    msg_ok2 = "Ditt lösenord har ändrats till: ",
    msg_min_length = "Lösenordet måste innehålla minst %s tecken",
    msg_max_length = "Lösenordet får maximalt innehålla %s tecken",

    help_title = "cmd_setpass.lua",
    help_usage = "[+!#]setpass nick <ANVÄNDARNAMN> <LÖSENORD>  /  [+!#]setpass nick myself <LÖSENORD>",
    help_desc = "Anger lösenord på en användare eller på dig själv",

    ucmd_menu_ct1_0 = { "Användare", "Kontroll", "Ändra", "Lösenord", "efter ANVÄNDARNAMN" },
    ucmd_menu_ct1_1 = { "Om dig", "ändra Lösenord" },
    ucmd_menu_ct1_2 = "Användare",
    ucmd_menu_ct1_3 = "Kontroll",
    ucmd_menu_ct1_4 = "Ändra",
    ucmd_menu_ct1_5 = "Lösenord",
    ucmd_menu_ct1_6 = "efter Användarnamn från lista",
    ucmd_menu_ct2_1 = { "Ändra", "Lösenord" },

    ucmd_pass = "Lösenord:",
    ucmd_nick = "Användarnamn:",

}