﻿return {

    help_title = "etc_topic.lua",
    help_usage = "[+!#]topic <NYTT-ÄMNE>|default",
    help_desc = "Anger nytt hubbämne eller återställer den till standard",

    msg_topic_changed = "%s har ändrat hubbämnet till: %s   |   det gamla hubbämnet var: %s",
    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_usage = "Användning: [+!#]topic <NYTT-ÄMNE>|default",
    msg_topic_reset = "%s  återställer hubbämnet till standard: %s",

    ucmd_popup = "Nytt ämne:",
    ucmd_menu = { "Hubb", "Kärna", "Hubbämne", "ändra ämne" },
    ucmd_menu2 = { "Hubb", "Kärna", "Hubbämne", "ändra till standard" },

}