﻿return {

    help_title = "cmd_myip.lua",
    help_usage = "[+!#]myip [<ANVÄNDARNAMN>]",
    help_desc = "Visar IP-adressen på en användare eller på dig själv",

    ucmd_menu_ct1 = { "Om dig", "visa IP" },
    ucmd_menu_ct2 = { "Visa", "IP" },

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_ip = "Din IP-adress är: ",
    msg_targetip = "Användarnamn: %s  |  IP: %s",

}