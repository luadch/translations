﻿return {

    block_msg = "Du har blivit bannad i %s minuter därför att du har DHT aktiverad i din klient. Inaktivera DHT och anslut igen när bann-tiden löpt ut.",
    report_msg = "%s blev bannad i %s minuter därför att DHT var aktiverat.",

}