﻿return {

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_userlist = "Användarlista:",
    msg_useramount = "Användare i varje åtkomstnivå:\n",

    help_title = "cmd_userlist.lua",
    help_usage = "[+!#]userlist [bydate]",
    help_desc = "Visar en lista över registrerade användare",


    ucmd_menu = { "Hubb", "etc", "Användarlista", "efter ÅTKOMSTNIVÅ" },
    ucmd_menu_bydate = { "Hubb", "etc", "Användarlista", "efter DATUM" },

}