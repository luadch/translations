﻿return {

    msg_invalid = "Ogiltigt hubbantal.",
    msg_max = [[


=== HUBBKONTROLL FÖR ANVÄNDAREN ===================

Du har blivit frånkopplad därför att:

Tillåtna publika hubbar: %s  |  du är i: %s
Tillåtna registrerade hubbar: %s  |  du är i: %s
Tillåtna operatörshubbar: %s  |  du är i: %s

Maximalt tillåtna hubbar: %s  |  du är i: %s

=================== HUBBKONTROLL FÖR ANVÄNDAREN ===
  ]],

    report_msg = "%s blev bannad i %s minuter därför att hubbegränsningen har överskridits. Hubbar: %s",
    msg_reason = "Överskrider hubbens användarantal",

}