﻿return {

    help_title = "cmd_reload.lua",
    help_usage = "[+!#]reload",
    help_desc = "Laddar om konfigurationen: cfg.tbl, user.tbl och alla skript",

    ucmd_menu = { "Hubb", "Kärna", "Ladda om hubben" },

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_ok = "Konfigurationen är omladdad.",

}