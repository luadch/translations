﻿return {

    help_title = "cmd_restart.lua",
    help_usage = "[+!#]restart",
    help_desc = "Startar om hubben",

    ucmd_menu = { "Hubb", "Kärna", "Hubbomstart", "KLICK" },

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_ok = "Hubben är omstartad.",
    
    msg_countdown = "*** Omstart av hubben om ***",

}