﻿return {

    help_title = "usr_hide_share.lua",
    help_usage = "[+!#]hideshare <ANVÄNDARNAMN>",
    help_desc = "Göm/visa utdelningen för en användare",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_isbot = "Användaren är en bot.",
    msg_notonline = "Användaren är frånkopplad.",
    msg_usage = "Användning: [+!#]hideshare <ANVÄNDARNAMN>",

    msg_default = "Åtkomstnivån bestämmer att denna användares utdelning är gömd.",
    msg_hide_user = "Utdelning är gömd för: %s",
    msg_hide_target = "Din utdelning gömdes av: %s",
    msg_unhide_user = "Utdelningen visas igen för: %s  |  Användaren blev frånkopplad",
    msg_unhide_target = "Din utdelning har återställts av: %s  |  Därför kommer du att bli frånkopplad nu",

    ucmd_menu_ct2_1 = { "Ändra", "Utdelning", "göm//visa igen" },

}