﻿return {

    help_title = "cmd_uptime.lua",
    help_usage = "[+!#]uptime",
    help_desc = "Visar din och hubbens drifttid",
    
    msg_denied = "Du har inte behörighet att använda detta kommando.",

    msg_years = " år, ",
    msg_days = " dagar, ",
    msg_hours = " timmar, ",
    msg_minutes = " min, ",
    msg_seconds = " sek",
    
    msg_unknown = "<OKÄNT>",
    
    msg_uptime = [[

    
=== DRIFTTID ==========================================================

                  Hubbens drifttid (sammanlagt):  %s
                  Hubbens drifttid (sen omstart):  %s
                  
                  Din drifttid:  %s

========================================================== DRIFTTID ===
  ]],

}