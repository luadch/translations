﻿return {

    help_title = "cmd_talk.lua",
    help_usage = "[+!#]talk <MEDDELANDE>",
    help_desc = "Prata i huvudchatten utan användarnamn",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    ucmd_menu = { "Användare", "Meddelande", "Prata" },
    ucmd_what = "Meddelande:",

}