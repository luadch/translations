﻿return {

    msg_invalid = "Ogiltigt hubbantal.",
    msg_max = [[

=== HUBBKONTROLL FÖR ANVÄNDAREN ===================

Du har blivit frånkopplad därför att:

Tillåtna publika hubbar: %s  |  du är i: %s
Tillåtna registrerade hubbar: %s  |  du är i: %s
Tillåtna operatörshubbar: %s  |  du är i: %s

Maximalt tillåtna hubbar: %s  |  du är i: %s

=================== HUBBKONTROLL FÖR ANVÄNDAREN ===
  ]],

    block_msg = "Du har blivit bannad i %s minuter därför att du överskridit hubbegränsningen. Kontrollera detta och försök igen när bann-tiden löpt ut.",
    report_msg = "%s blev bannad i %s minuter därför att hubbegränsningen har överskridits.",

}