﻿return {

    help_title = "usr_redirect.lua",
    help_usage = "[+!#]redirect <ANVÄNDARNAMN> <URL>",
    help_desc = "Omdirigera användare till URL",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_usage = "Användning: [+!#]redirect <ANVÄNDARNAMN> <URL>",
    msg_god = "Du har inte behörighet att omdirigera denna användaren.",
    msg_isbot = "Användaren är en bot.",
    msg_notonline = "Användaren är frånkopplad.",
    msg_redirect = "[ OMDIRIGERA ]--> Användaren:  %s  |  har omdirigerats till:  %s",
    msg_report_redirect = "[ OMDIRIGERA ]--> Användaren:  %s  |  har omdirigerat användaren:  %s  |  till:  %s",

    ucmd_menu_ct2_1 = { "Omdirigera", "standard URL" },
    ucmd_menu_ct2_2 = { "Omdirigera", "egen URL" },
    ucmd_url = "URL för omdirigering:",

    msg_report = "[ OMDIRIGERA ]--> Användaren:  %s  |  med åtkomstnivå  %s [ %s ]  |  har automatiskt omdirigerats till:  %s",

}