return {

    warning = [[


=== VARNING ============================================================

               Standard hubbägarkontot 'dummy' är fortfarande aktiverat! Inaktivera det så fort som möjligt!

============================================================ VARNING ===
  ]],

}