﻿return {

    msg_denied = "Du har inte behörighet att använda detta kommando eller att ta bort användarkonton med denna åtkomstnivå.",
    msg_import = "Ett fel uppstog vid importering av tilläggsmodul.",
    msg_usage = "Användning: [+!#]delreg nick <ANVÄNDARNAMN>  /  eller radera med svartlistspost:  [+!#]delreg nick <ANVÄNDARNAMN> <BESKRIVNING>",
    msg_error = "Ett fel uppstod: ",
    msg_del = "Ditt konto är raderat.",
    msg_bot = "Fel: Användaren är en bot.",
    msg_ok = "Användaren  %s  har blivit raderad av  %s",
    msg_ok2 = "%s  blev raderad och svartlistad av  %s  anledning: %s",
    msg_notfound = "Användaren är inte registrerad.",

    help_title = "cmd_delreg.lua",
    help_usage = "[+!#]delreg nick <ANVÄNDARNAMN>  /  eller radera med svartlistspost:  [+!#]delreg nick <ANVÄNDARNAMN> <BESKRIVNING>",
    help_desc = "Raderar en användare",

    ucmd_menu_ct1 = { "Användare", "Kontroll", "Delreg", "efter ANVÄNDARNAMN" },
    ucmd_menu_ct2 = { "Delreg", "OK" },
    ucmd_nick = "Användarnamn:",
    ucmd_reason = "Anledning: (läggs inte i svartlistan om den är tom)",

}