﻿return {

    report_msg = "%s blev bannad i %s minuter därför att DHT var aktiverat.",
    msg_reason = "DHT är aktivt",

}