﻿return {

    msg_motd = [[


=== MOTD ========================================================================================

                                                                     Välkommen %s
                                                                     Detta är dagens information (MOTD)

======================================================================================== MOTD ===
      ]], -- det går att lägga till %s för att få med användarnamnet i texten

}