﻿return {

    msg_slotlimits = "Minsta antal slots: %s  |  Max antal slots: %s  |  Dina slots: %s",

}