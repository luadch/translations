﻿return {

    msg_denied = "Du har inte behörighet använda detta kommando.",
    msg_import = "Ett fel uppstog vid importering av tilläggsmodul.",
    msg_report = "Användaren %s registrerade %s med åtkomstnivå %d [ %s ]",
    msg_level = "Du har inte behörighet att registrera på denna åtkomstnivå.",
    msg_usage = "Användning: +reg nick <ANVÄNDARNAMN> <ÅTKOMSTNIVÅ>",
    msg_error = "Ett fel uppstod: ",
    msg_ok = "Användare registrerades med följande  parametrar: Användarnamn: %s | Lösenord: %s | Åtkomstnivå: %s [ %s ]",
    msg_accinfo = [[


=== KONTO ========================================

    Användarnamn: %s
    Lösenord: %s

    Åtkomstnivå: %s  [ %s ]
    
    Hubbnamn: %s
    Hubbadress: %s
    
======================================== KONTO ===

        ]],

    help_title = "cmd_reg.lua",
    help_usage = "[+!#]reg nick <ANVÄNDARNAMN> <ÅTKOMSTNIVÅ>",
    help_desc = "Registrera en ny användare",

    ucmd_menu_ct1_1 = "Användare",
    ucmd_menu_ct1_2 = "Kontroll",
    ucmd_menu_ct1_3 = "Registrera",
    ucmd_menu_ct2 = { "Registrera", "OK" },
    ucmd_passwort = "Lösenord:",
    ucmd_level = "Åtkomstnivå:",
    ucmd_nick = "Användarnamn:",
    
    msg_blacklist1 = "Fel: Denna användaren är svartlistad!",
    msg_blacklist2 = "Anledning: ",
    msg_blacklist3 = "Borttagen på: ",
    msg_blacklist4 = "Borttagen av: ",

}