﻿return {

    msg_usage = "Användning:",
    msg_description = "Beskrivning:",
    msg_minlevel = "Lägsta åtkomstnivå:",

    help_title = "cmd_help.lua",
    help_usage = "[+!#]help",
    help_desc = "Visa denna hjälp för hubbkommandon",

    ucmd_menu = { "Allmänt", "Hjälp" },
    
    msg_out = [[


=== TILLGÄNGLIGA KOMMANDON =================================================================================
%s
================================================================================= TILLGÄNGLIGA KOMMANDON ===
  ]],

}